module parser